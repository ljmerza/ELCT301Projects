opamp circuit
.lib eval.lib

X1 0 2 4 5 3 LM324
VS 1 0 PULSE(0 1 0 10nS 10nS .8e-3 1.6e-3) Ac 1
* V3 1 0 AC 1
R1 1 2 1K 
RF 2 3 10K
V1 4 0 15V
V2 5 0 -15V

.AC DEC 100 1Hz 1MEG
.PROBE
.END

