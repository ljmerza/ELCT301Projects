Diode Current Source
.lib eval.lib

VCC 1 0 15V
R1 1 2 20k
RL 1 3 10k
Q1 3 2 0 Q2N2222
Q2 2 2 0 Q2N2222
.MODEL Q2N2222 NPN(BF=300)

.TRAN 10us 2ms
.PROBE
.END