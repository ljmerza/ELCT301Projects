Bouncing Switch
* File bounceswitch.cir

S1 1 0 2 0 SMOD


.MODEL SMOD VSWITCH(RON=1)

R1 3 1 1K
VCC 3 0 DC 5V
V2 4 0 PWL(1E-3 0V 1.0001E-3 5V 1.01E-3 5V 1.0101E-3 0V 1.02E-3 0V 1.0201E-3 5V 1.03E-3 5V 1.0301E-3 0V 1.04E-3 0V 1.0401E-3 5V )

V3 2 4 PWL(2E-3 0V 2.0001E-3 -5V 2.01E-3 -5V 2.0101E-3 0V 2.02E-3 0V 2.0201E-3 -5V 2.03E-3 -5V 2.0301E-3 0V 
+    2.04E-3 0V 2.0401E-3 -5V )


.TRAN 20E-6 3E-3 
.PROBE
.END
