One Transistor Current Source
.lib eval.lib

VCC 1 0 15V
RL 1 3 10k
R1 1 2 2.35Meg
Q1 3 2 0 Q2N2222
.MODEL Q2N2222 NPN(BF=300)

.TRAN 10us 2ms
.PROBE
.END