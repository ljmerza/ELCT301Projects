signal generator at 10Hz
.LIB eval.lib
VCC 15 0 15V
VEE 16 0 -15V

*Schmitt Trigger
R300 1 2 100k
R301 2 4 100k
X1 2 0 15 16 3 LM324
R302 3 4 1k
D300 5 4 D1N750 
D302 5 0 D1N750 
*set to operate at 10 Hz
R310 4 6 1k
RFREQ 6 7 249k
*comment out above two lines and uncomment following line to operate at 2500 Hz
*R310 4 7 1k

*Integrator
X2 0 7 15 16 8 LM324
C310 7 8 100n IC=5V
R320 8 9 3.3k
R321 9 0 1.8k
RJUMP300 1 8 100
X3 9 10 15 16 10 LM324

*Diode wave shaping circuit
R330 10 11 1k
D330 12 11 D1N4148 
D331 11 12 D1N4148 
R331 12 0 2.7k
D332 13 11 D1N4148 
D333 0 13 D1N4148 
D334 11 14 D1N4148 
D335 14 0 D1N4148

.TRAN 5ns .2s
.FOUR 10Hz V(11)
.PROBE
.END
