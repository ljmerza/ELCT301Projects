555d Astable Simulation
.lib eval.lib

Vcc 1 0 DC 5V

R1 1 3 100K
R2 3 4 10K
RL 5 0 1K

C1 4 0 47uF
C2 2 0 10nF

X1 0 4 5 1 2 4 3 1 555d

.TRAN 1e-3 20  
.PROBE
.END
