555d Monostable Simulation
.lib eval.lib

Vcc 1 0 DC 5V
Vi 5 0 PULSE(5 0 5ms 1us 1us 1ms 10ms)

R1 1 2 500K
RL 4 0 1K
C1 2 0 10nF
C2 3 0 10nF

X1 0 5 4 1 3 2 2 1 555d

.TRAN 1ms 40ms  
.PROBE
.END
